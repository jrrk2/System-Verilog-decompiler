
module test_initial(
  output logic q
);
  initial
    q = 1'b0;
endmodule
